a     a   v     <  �  �    7  _  t  }  �  �  �  �      (  �  �  �  �     v   FileAndType�     �{"baseDir":"/home/alex/Repos/Harvest-Grove/Documentation","file":"api/City.NPC.NPCDialogueUI.yml","type":"article","sourceDir":"api/","destinationDir":"api/"}   <  OriginalFileAndType�   �  �{"baseDir":"/home/alex/Repos/Harvest-Grove/Documentation","file":"api/City.NPC.NPCDialogueUI.yml","type":"article","sourceDir":"api/","destinationDir":"api/"}   �  Key*      ~/api/City.NPC.NPCDialogueUI.yml   7  LocalPathFromRoot(   _  api/City.NPC.NPCDialogueUI.yml   t  LinkToFiles	   }     �  
LinkToUids=   �  �    .  o  �  �  �    !  C  n  �  �  I     ?City.NPC.NPCDialogueUI.Construct(ICanvasData,IInventoryService)   .  System.ObjectA   o  7City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button@)9   �  /City.NPC.NPCDialogueUI.InstantiateChoiceButton*   �  Global.ICanvasData+   �  !City.NPC.NPCDialogueUI.CloseNpcUI     City.NPC    !  City.NPC.NPCDialogueUI"   C  Global.IInventoryService+   n  !City.NPC.NPCDialogueUI.Construct*,   �  "City.NPC.NPCDialogueUI.CloseNpcUI*    �  Global.TextMeshProUGUI   �  Global.Button   �  FileLinkSources   �  {}     UidLinkSources     {}   (  Uids�  �  �[{"name":"City.NPC.NPCDialogueUI","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.Construct(ICanvasData,IInventoryService)","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button@)","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.CloseNpcUI","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.Construct*","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.InstantiateChoiceButton*","file":"api/City.NPC.NPCDialogueUI.yml"},{"name":"City.NPC.NPCDialogueUI.CloseNpcUI*","file":"api/City.NPC.NPCDialogueUI.yml"}]   �  ManifestProperties   �  {}   �  DocumentType	      ^0  d8  {"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.PageViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","items":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"City.NPC.NPCDialogueUI","commentId":"T:City.NPC.NPCDialogueUI","id":"NPCDialogueUI","isEii":false,"isExtensionMethod":false,"parent":"City.NPC","children":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["City.NPC.NPCDialogueUI.CloseNpcUI","City.NPC.NPCDialogueUI.Construct(ICanvasData,IInventoryService)","City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button@)"]},"langs":{"$type":"System.String[], System.Private.CoreLib","$values":["csharp","vb"]},"name":"NPCDialogueUI","nameWithType":"NPCDialogueUI","fullName":"City.NPC.NPCDialogueUI","type":"Class","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"NPCDialogueUI","path":"","startLine":8879,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["cs.temp.dll"]},"namespace":"City.NPC","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public class NPCDialogueUI : MonoBehaviour","content.vb":"Public Class NPCDialogueUI Inherits MonoBehaviour"},"inheritance":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["System.Object"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"City.NPC.NPCDialogueUI.Construct(ICanvasData,IInventoryService)","commentId":"M:City.NPC.NPCDialogueUI.Construct(ICanvasData,IInventoryService)","id":"Construct(ICanvasData,IInventoryService)","isEii":false,"isExtensionMethod":false,"parent":"City.NPC.NPCDialogueUI","langs":{"$type":"System.String[], System.Private.CoreLib","$values":["csharp","vb"]},"name":"Construct(ICanvasData, IInventoryService)","nameWithType":"NPCDialogueUI.Construct(ICanvasData, IInventoryService)","fullName":"City.NPC.NPCDialogueUI.Construct(ICanvasData, IInventoryService)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"Construct","path":"","startLine":8910,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["cs.temp.dll"]},"namespace":"City.NPC","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public void Construct(ICanvasData canvas, IInventoryService inventoryService)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"canvas","type":"Global.ICanvasData"},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"inventoryService","type":"Global.IInventoryService"}]},"content.vb":"Public Sub Construct(canvas As ICanvasData, inventoryService As IInventoryService)"},"overload":"City.NPC.NPCDialogueUI.Construct*"},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button@)","commentId":"M:City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button@)","id":"InstantiateChoiceButton(Button@)","isEii":false,"isExtensionMethod":false,"parent":"City.NPC.NPCDialogueUI","langs":{"$type":"System.String[], System.Private.CoreLib","$values":["csharp","vb"]},"name":"InstantiateChoiceButton(out Button)","nameWithType":"NPCDialogueUI.InstantiateChoiceButton(out Button)","fullName":"City.NPC.NPCDialogueUI.InstantiateChoiceButton(out Button)","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"InstantiateChoiceButton","path":"","startLine":9163,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["cs.temp.dll"]},"namespace":"City.NPC","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"protected TextMeshProUGUI InstantiateChoiceButton(out Button choiceBtnButton)","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","id":"choiceBtnButton","type":"Global.Button"}]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"Global.TextMeshProUGUI"},"content.vb":"Protected Function InstantiateChoiceButton(choiceBtnButton As Button) As TextMeshProUGUI"},"overload":"City.NPC.NPCDialogueUI.InstantiateChoiceButton*","nameWithType.vb":"NPCDialogueUI.InstantiateChoiceButton(Button)","fullName.vb":"City.NPC.NPCDialogueUI.InstantiateChoiceButton(Button)","name.vb":"InstantiateChoiceButton(Button)"},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"City.NPC.NPCDialogueUI.CloseNpcUI","commentId":"M:City.NPC.NPCDialogueUI.CloseNpcUI","id":"CloseNpcUI","isEii":false,"isExtensionMethod":false,"parent":"City.NPC.NPCDialogueUI","langs":{"$type":"System.String[], System.Private.CoreLib","$values":["csharp","vb"]},"name":"CloseNpcUI()","nameWithType":"NPCDialogueUI.CloseNpcUI()","fullName":"City.NPC.NPCDialogueUI.CloseNpcUI()","type":"Method","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","id":"CloseNpcUI","path":"","startLine":9265,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":["cs.temp.dll"]},"namespace":"City.NPC","summary":"<p sourcefile=\"api/City.NPC.NPCDialogueUI.yml\" sourcestartlinenumber=\"2\">Closes the NPC panel UI</p>\n","example":{"$type":"System.Collections.Generic.List`1[[System.String, System.Private.CoreLib]], System.Private.CoreLib","$values":[]},"syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public void CloseNpcUI()","content.vb":"Public Sub CloseNpcUI()"},"overload":"City.NPC.NPCDialogueUI.CloseNpcUI*"}]},"references":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC","commentId":"N:City.NPC","name":"City.NPC","nameWithType":"City.NPC","fullName":"City.NPC","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City","name":"City","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":".","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC","name":"NPC","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], System.Private.CoreLib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City","name":"City","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":".","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC","name":"NPC","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","commentId":"T:System.Object","parent":"System","isExternal":true,"name":"object","nameWithType":"object","fullName":"object","nameWithType.vb":"Object","fullName.vb":"Object","name.vb":"Object"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System","commentId":"N:System","isExternal":true,"name":"System","nameWithType":"System","fullName":"System"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC.NPCDialogueUI.Construct*","commentId":"Overload:City.NPC.NPCDialogueUI.Construct","name":"Construct","nameWithType":"NPCDialogueUI.Construct","fullName":"City.NPC.NPCDialogueUI.Construct"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"Global.ICanvasData","isExternal":true,"name":"ICanvasData","nameWithType":"ICanvasData","fullName":"ICanvasData"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"Global.IInventoryService","isExternal":true,"name":"IInventoryService","nameWithType":"IInventoryService","fullName":"IInventoryService"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC.NPCDialogueUI.InstantiateChoiceButton*","commentId":"Overload:City.NPC.NPCDialogueUI.InstantiateChoiceButton","name":"InstantiateChoiceButton","nameWithType":"NPCDialogueUI.InstantiateChoiceButton","fullName":"City.NPC.NPCDialogueUI.InstantiateChoiceButton"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"Global.Button","isExternal":true,"name":"Button","nameWithType":"Button","fullName":"Button"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"Global.TextMeshProUGUI","isExternal":true,"name":"TextMeshProUGUI","nameWithType":"TextMeshProUGUI","fullName":"TextMeshProUGUI"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"City.NPC.NPCDialogueUI.CloseNpcUI*","commentId":"Overload:City.NPC.NPCDialogueUI.CloseNpcUI","name":"CloseNpcUI","nameWithType":"NPCDialogueUI.CloseNpcUI","fullName":"City.NPC.NPCDialogueUI.CloseNpcUI"}]},"shouldSkipMarkup":false,"_appFooter":"Harvest Grove ","_appTitle":"Harvest Grove code documentation","_enableSearch":true,"_systemKeys":{"$type":"System.String[], System.Private.CoreLib","$values":["uid","isEii","isExtensionMethod","parent","children","href","langs","name","nameWithType","fullName","type","source","documentation","assemblies","namespace","summary","remarks","example","syntax","overridden","overload","exceptions","seealso","see","inheritance","derivedClasses","level","implements","inheritedMembers","extensionMethods","conceptual","platform","attributes","additionalNotes"]}}�   	9  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, System.Private.CoreLib],[System.Object, System.Private.CoreLib]], System.Private.CoreLib"}	   9   